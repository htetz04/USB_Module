`timescale 1ns/10ps


module USB_TX_Packet_Loader(

);

endmodule